class ahb_tx extends uvm_sequence_item;
  rand bit [31:0] addr;
  rand bit [31:0] addr_t;
  rand bit [31:0] dataQ[$];
  rand bit wr_rd;
  //rand bit [2:0] burst;
  rand burst_t burst;
  rand bit [2:0] size;
  rand bit [4:0] len;
  rand bit [6:0] prot;
  rand bit excl;
  rand bit [3:0] master;
  rabd bit nonsec;
  rand bit mastlock;
  bit [1:0] resp;
  bit exokay;
  
  integer txsize;
  bit [31:0] lower_wrap_addr;
  bit [31:0] upper_wrap_addr;
  
  // htrans, hready & hreadyout are handshaking signals
  // herror is generated by slave
  // no clk and rst as well (hclk and hrst)
  // leaving h out makes it generic for other protocols
  
  `uvm_object_utils_begin(ahb_tx)
  `uvm_field_int(addr, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_queue(dataQ, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_int(wr_rd, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_enum(burst_t, burst, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_int(size, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_int(len, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_int(prot, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_int(excl, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_int(master, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_int(nonsec, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_int(mastlock, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_int(resp, UVM_ALL_ON | UVM_NOPACK)
  `uvm_field_int(exokay, UVM_ALL_ON | UVM_NOPACK)
  `uvm_object_utils_end
  
  `NEW_OBJ
  
  function void post_randomize();
    addr_t = addr;
    calc_wrap_boundaries();
  endfunction
  
  //Constraints
  
  constraint burst_len_c {
    (burst == SINGLE) -> (len == 1);
    (burst inside {INCR4, WRAP4} -> (len == 4);
    (burst inside {INCR8, WRAP8} -> (len == 8);
    (burst inside {INCR16, WRAP16} -> (len == 16);
     len inside {[1:16]}; //taking care of INCR burst
  }
  
  constraint dataQ_c {
    dataQ.size() == len;
  }
     
  //AHB only supports aligned transfers
  constraint aligned_c {
    addr % (2**size) == 0;
  }
  
  //keep default transfers as INCR4
  constraint burst_c {
    soft burst == INCR4; //if user doesn't give any specific constraint for burst then use this default value
  }
     
  constraint size_c {
    soft size == 2; //4 bytes per beat => fit into 32 bit data bus
  }
  
  constraint master_c {
    soft master == 0;  
  }
     
  //Methods
  //wrap boundaries
     
  function void calc_wrap_boundaries();
    //txsize = num_transfers(beats) * bytes_per_beat;
    txsize = len * (2**size); //wrap boundaries will be 0, 1*txsize, 2*txsize...
    //0, 64, 128
    //78 => 78
    lower_wrap_addr = addr - (addr%txsize);
    	//78 - 78%64 = 78 - 14 = 64
    upper_wrap_addr = lower_wrap_addr - txsize - 1;
    	//64 + 64 - 1 = 127
  endfunction
  
endclass
     

/*General Transaction class:
1) properties (fields required to implement all the aspects of (AHB) transactions)
2) methods
	. copy, print, compare => these methods come due to automatic registration of fields into the factory
	. pack, unpack? NO
		. AHB is not a serial protocol
		. only serial protocols require PACK, UNPACK     methods
	. what other methods are required?
		. method for calculating wrap boundaries for given address
3) constraints

I declared all the fields of the AHB interface except for the handshaking signals, clk and rst signals

handshaking signals: htrans, hready and hreadyout
clock & reset: hclk, hrst

resp, exokay are non rand because these are driven by the slave. Any signals driven by the slave can't be declared as rand.

Coding transaction class efficiently is important for any testbench development, so that you can cover all features properly, and can implemented transaction related methods properly (instead of implementing elsewhere) as well as constraints. It makes tb dev easier.

You can code way more constraints and methods.